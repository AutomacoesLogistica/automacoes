��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  9yS�    GND      �  9YJg    5V      �  �q�    12V / 5V      �  �Y�g    LM2596      �  �a~o    MIKE(2) - 1=12v   -   2 = GND      �  Aq�    Entrada 12V      �  9hG    MIKE(4) - Pino4      �  � h    MIKE(4) - Pino3      �  i ���    :MIKE(8) - 1_12V(Marrom)  - 2_Sinal(Preto) - 3 GND ( Azul )      �  � 18?    MIKE(4) - Pino1      �  � �8�    MIKE(4) - Pino2      �  ��y�    &GPIO saida para pulso abertura cancela      �  ��'    Pulso para abrir cancela ( 12 )      �  I�W    'Sinal pulso cancela vindo do totem (13)      �  �&�    :Sinal entrada sensor vandalismo da cancela ESP32 Lora (23)      �  �     7Sinal entrada Aberta/Fechado da cancela ESP32 Lora (17)      �   a� o    *Rele sinal de pulso cancela vindo do totem      �  � �=�    Representando sensor vandalismo      �  � 	`    ,Rele sinal entrada Aberta/Fechado da cancela                    ��� 	 CRailThru�� 	 CTerminal  �-�     0 d                   �  �1�     4                       |.�         ����    ��  h-i     0 d                   �  h1i     3                       d.l     "    ����    ��  ����     1 d                   �  ����     2                       �|��     %    ����    ��  �h�i     / d                   �  �h�i     2                       �d�l     (    ����    ��  x	�      0 d                   �  |	�     -                       z�    +    ����    ��  P	e      + d        �          �  T	i     0                       Rf    .    ����    ��  �x��      2 d                   �  �|��     .                       �z��    1    ����    ��  �P�e      , d                   �  �T�i     2                       �R�f    4    ����    ��  ����     . d                   �  ����     -                       ����     7    ����    ��  �P�Q     , d                   �  �P�Q     +          �            �L�T     :    ����    ��  CBattery��  CValue  #�K�    3.3V(    ffffff
@      �? V �  XhY}      %   ffffff
@%�]���  �  X�Y�     !           %�]��>    L|d�     @    ��      ��  �        d        �          �  �      *                       ��      C    ����    ��  �@A     # d        �          �  �@A     )                       �<D     F    ����    ��  ����     ( d n�ݑYH�?          �  ����     '   n�ݑYH�?            ����     I    ����    ��  CEarth�  ����      ! 	            �OU<    ����     M    ��      �� 	 CResistor>�  �v��    1k        @�@      �?k  �  ����     &   n�ݑYH�?          �  p���     '   n�ݑYH�?            ����    Q    ��      ��  CNPN��  CDummyValue  �x�x    100hFE            Y@      �? hFE �  �h�}      " 	 AQRff
@z�_��>  �  ����     & 	 n�ݑYH�?    TY�;  �  ����     !           �  _���    �|��     W    ��      ��  CDiode�  �h�i     "   AQRff
@�|�Q��  �  �h�i     %   ffffff
@�|�Q�=    �\�t    \    ��      �� 
 CRelaySPDT�  �8�9                �          �  �P�Q     %   ffffff
@B|iP��>  �  �P�Q     "   AQRff
@B|iP���  �  �@�A     #          �          �  �0�1     $                       �,�X    `    ��      K��  ����                 �Q9�2F>    ����     f    ��      K��  0�1�       	                     #�;�     h    ��      N�>�  @�`�    1k        @�@      �?k  �  \�q�               �          �  0�E�                            D�\�    k    ��      �� 	 CVoltRail>�   �C �    12V(          (@      �? V �  L �a �             (@            D �L �     p    ����     ^��  ` �u �      	       (@          �  ` �u �       �,   "@�9�NۻS�  �  � �� �       �,   "@�9�NۻS<  �  � �� �               �          �  � �� �             (@            t �� �    r    ��      <�>�   �3 �    9V(          "@      �? V �  @ �A �        �,   "@�9�NۻS<  �  @ �A �      	 [8Z6>rO�8l�>�    4 �L �     y    ��      Z��  � �� �       �,   "@          �  ` �u �       �,   "@            t �� �    |    ��      ��  CSPST��  CToggle  P �p          �  @ �U �        [8Z6>          �  l �� �       �,   "@            T �l �     �      ��    K��  h�i�       	                     [�s�     �    ��      �� 
 CVoltmeter��  CMeter  3�[�     3.30(    �  hxi�         ���df
@          �  h�i�                            \�t�     �    ��      K��  `a       	                     Sk$     �    ��      ����  +�S�     3.30(    �  `�a�         ���df
@          �  `�a	                            T�l�     �    ��      m�>�  + � S �     12V(          (@      �? V �  \ � q �              (@            T � \ �      �    ����     ~���  8 �X �     �   �  ( �= �                ��J=
��  �  T �i �                ��J=
�?    < �T �     �     ��    Z��  t x� y                r��{���  �  H x] y             "@r��{��=    \ lt �    �    ��      <�>�  ��y �    9V(          "@      �? V �  ( `) u              "@��J=
��  �  ( �) �      	         ��J=
�?     t4 �     �    ��      ^��  H H] I             (@          �  H `] a             "@
8\=
�?  �  t `� a                
8\=
��  �  t P� Q             (@          �  t @� A               �            \ <t h    �   ��      ����  #9KG     3.30(    �  X Y5      
   ���df
@          �  XLYa                            L4dL     �    ��      K��  X`Yu       	                     Ktc|     �    ��      N�>�  ��,    1k        @�@      �?k  �  �0�1        ffffff
@�ʡ寘->  �  �0�1     
   ���df
@�ʡ寘-�    �,�4    �    ��      N�>�  ���    1k        @�@      �?k  �  ��	        ffffff
@�ʡ寘->  �  ��	        ���df
@�ʡ寘-�    ��    �    ��      N�>�  �f�t    1k        @�@      �?k  �  �x�y        ffffff
@�ʡ寘->  �  �x�y        ���df
@�ʡ寘-�    �t�|    �    ��      K��   X!m      	 	                     l+t     �    ��      N�>�  0FPT    1k        @�@      �?k  �  LXaY               �          �   X5Y     	                       4TL\    �    ��      m�>�  � �     9V(          "@      �? V �  � � 	             "@            � �      �    ����     �� 	 CIsolator�  �x��         ���df
@e¡寘->  �  pxq�                �          �  p�q�      	        �          �  ����                e¡寘-�    d���     �    ��      ��  CFloatSwitch��  CWaterLevel  � 0    	 �   �  � � 	      	       "@          �  !	               �            �      �     ��    ���  ��         ���df
@e¡寘->  �  pq                �          �  p4qI               �          �  �4�I                e¡寘-�    d�4     �    ��      m�>�  C� k�     3.3V(    ffffff
@      �? V �  t� ��         ffffff
@X9�2F�    l� t�      �    ����     K��  h	}                             � |�     �    ��      N�>�  8nX|    1k        @�@      �?k  �  T�i�               �          �  (�=�                            <|T�    �    ��      ���  �0�E      
   ���df
@e¡寘->  �  h0iE                �          �  h\iq               �          �  �\�q                e¡寘-�    \D�\     �    ��                    ���  CWire  x�      0 �  xy     0 ��� 
 CCrossOver  ����        �0�	       �  hi     0 �  �x�y     2 �  �x��      2 �  ����     2 �  �h�y      2 �  �h�i     2 �  ��1      
 �  ����     . �  �P�Q     , �  �P	Q     + �  h	y      0 �  ��	�     - ��  ��        �Y     
 �  � @QA      �  � �Q�      ��  n�t�        X���     ! ��  n�t�        p�q�      ' �  Xh�i     % �  � �       �  � �9        �  �@�A     # �  ��q�     ' �  �P�i      " �  �P�i      % �  Pxqy      �  PxQ�       ��  �t�|      �  �\�d        �H��       ��  ����      �  ��        �p�I       �  �H�I      �  ����      �  �p�q      ��  �t�|        �x�y      ��  �\�d      �  �\�d        �`ia      ��  ��        ��	      ��  ����      �  ����        ��a�      �  h`iy       �  �`�y       ��  �\�d        ��y       �  ` �a �       �  @ �a �      �  � �� �       �  � �� �       �  � �� �      �  ���	       �  P0i1      �  P0QA       �  hpi�       �  H (I I       �  H (q )      �  p � q )       �  h �� �      �  � x� �       �  � `� y       �  ( `I a      �  H `I y       �  XY!      
 ��  ��        �� �1       �  �� ��       �  �0�1     
 �   q	      �  `XqY      �  pHqY       �  (h)�       �  h)i                    �                            �        � " # #     % & & �   ( ) ) � � + , , � � . / / � � 1 2 2 � � 4 5 5 � � 7 8 8 � � : ; ; � @ � @ A A � � C D D   � F G G     I J J � M Y M Q Q X R � R W \ W X Q X Y Y � \ \  ] ] ` � ` a a b b  c c � d d   f f h l h k k � l h l p p r r p r s s t t u u � v v   y y z z � | | } } � z � � � � � � � � � � � � � � � � � � � � � &� � � � � '� � )� +� � *� � � � � $� � +� � � )� �   � � � � ,� � � � � � � � � -� 0� � � � � � � � � � � � � � � 2� � � � � � � � � � � � k � � � � � � � 1�  � � 1� � � 3� � 
� � /� 5� � � #� 4� � 0� � !� � � #� � �  � � � � � " � 1 � � & � � � ) 5 � � 2 7 4 : ; . / + 8 , � .� ,� "u � � A M � � R � @ ] � C � ` c F J � b W a � � � 
� � f � � 	� � �  � � � � � } y s t | � "� !� � � %� $&� %� (� '� (� � *� � � -� /� � -� � � � � 3� 25� � 4 5          �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 