��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  )I ^W     Mike(4) - 2      �  )� ^�     Mike(4) - 1      �  a � � �     Pino 5 - NC      �  a � � �     Pino 4 - Saida Corrente      �  a � � �     Pino 3 - GND      �  a � � �     Pino 2 - Saida Tensao      �  a � � �     Pino 1 - VCC 18 a 30V      �  Y�    
GPIO04 - 7      �  1ijw    
GPIO03 - 5      �  1� j�     
GPIO02 - 3      �  �i�w    Cooler      �  ����    5V      �  9�J�    5V      �  9y P�     3V3      �  �� �     Raspberry PI3 B+      �  )�R�    Pino 13      �  i9 �G     GND      �  	F    Mike(8) - 8      �  � F�     Mike(8) - 7      �  ����    Mike(8) - 3 e 4      �  Q���    Mike(8) - 1 e 2      �  	�P�    Mike(8) - 5 e 6      �  	�A�    	C - PRETO      �  ���    NA - VERMELHO      �  I���    
NF - VERDE      �  	Q>_    RELE 3V3      �  ����    
ESP32 LORA      �  y� ��     01DF100 IFM      �  iq �     24V                    ��� 	 CRailThru�� 	 CTerminal  h � } �       d        �          (�  l � � �                �            j � ~ �      )    ����    ��  CEarth(�  �	�                             ���     -    ��      &�(�  �H�I      d                   (�  �H�I                            �D�L     /    ����    &�(�  hHi]       d                   (�  hLia                            dJl^    2    ����    &�(�  hxi�       d                   (�  h|i�                            dzl�    5    ����    +�(�  ����                             ����     8    ��      &�(�  hP }Q       d                   (�  lP �Q                             jL ~T      :    ����    ��  CAND(�  P0 QE                 �          (�  @0 AE                 �          (�  H\ Iq                             <D T\     >      ��    &�(�  �       d                   (�  �                            �    B    ����    +�(�   ��                             ��     E    ��      &�(�  0�1�       d                   (�  0�1�                            ,�4�    G    ����    &�(�  0�1       d                   (�  0�1                            ,�4    J    ����    &�(�  ��       d                   (�  ��                            ��    M    ����    &�(�  (�)�       d                   (�  (�)�                            $�,�    P    ����    &�(�  @�A�       d                   (�  @�A�                            <�D�    S    ����    &�(�  H0IE       d                   (�  H4II                            D2LF    V    ����    &�(�  ����      d                   (�  ����                            �|��     Y    ����    &�(�  �� ��       d                   (�  �� ��                             �� ��      \    ����    +�(�  X�Y�                             K�c�     _    ��      &�(�  �� ��       d                   (�  �� ��                             �� ��      a    ����    &�(�  �� ��       d                   (�  �� ��                             �� ��      d    ����    &�(�   ��      d                   (�  ��     	                       ��     g    ����    &�(�  p���      d                   (�  t���                            r���     j    ����    +�(�  ����      
 	                     ���     m    ��      +�(�  � �5       	                     �4�<     o    ��      �� 	 CIsolator(�  ����                           (�  ����       	        �          (�  ����     
                     (�  ����     
                       ����     r    ��      �� 	 CResistor��  CValue  �i�w    10k          ��@      �?k  (�  �P�e                           (�  �|��                           �d�|     z    ��      v�x�  x���    100         Y@      �?   (�  ����               �          (�  h�}�     	                       |���    ~    ��      &�(�  h� }�       d                   (�  l� ��                             j� ~�      �    ����    &�(�  �� ��       d                   (�  �� ��                             �� ��      �    ����    &�(�  �� ��       d                   (�  �� ��                             �� ��      �    ����    &�(�  �� ��       d                   (�  �� ��                             �� ��      �    ����    &�(�  h� }�       d                   (�  l� ��                             j� ~�      �    ����    v�x�  x� ��     1k        @�@      �?k  (�  �� ��                �          (�  h� }�                             |� ��     �    ��      v�x�  �� ��     10k          ��@      �?k  (�  �� ��                            (�  �� ��                             �� ��      �    ��      p�(�  �� ��                            (�  �� ��        	        �          (�  ��!                          (�  ��!                            �� �     �    ��                    ���  CWire  � � 	�       ��  X � i �       ��  X � Y !       ��  X  	!      ��  � 	!       ��  @I      ��  0A      ��  @�A       ��  @���      ��  �p��       ��  hp�q      ��  h� iq       ��  hpi�       ��  ��	�      ��  ��      ��  `���      ��  �      ��  �	      ��  	I       ��  �H	I      ��  HI      ��  �H�I      ��  �H��       ��  H�       ���� 
 CCrossOver  �� ��         �P ��        ��  ����      ��  ���       ��  ���       ��  ��1�      ��  0�1�       ��  0�1�       ��  h`iy       ��  `�i�      ��  h�q�      ��  `�a�       ��  ���      ��  �� ��       ��  �P �Q       ��  ���      ��  H� i�       ��  �� I�       ��  Hp I�        ��  ��       ��   ��      ��         ��  1      ��  � �!      ��  ��1�      ��  0�Y�      ��  ����      ����  �� ��         �� i�       ��   ��      ��  �)�      ��  (�A�      ��  @�I�      ��  HHI�       ��   �       ��  HI1       ��  ����       ��  ����       ��  ����      ��  ����       ��  �� ��       ��  ����       ��  �� ��        ����  �� ��         �� ��       ��  �� ��        ��  �� ��        ��  �� ��        ����  �� ��         �� �Q       ��  X�i�      ��  �� ��        ��  �� ��       ��  �� ��        ��  �i�     	 ��   ��       ��   ��       ��  �� �       ��  �P�Q      ��  �� ��       ��  ����     
 ��  �� ��        ��  �� ��       ��  �� �!       ��  h� i�        ��  �� ��        ��  �� ��        ��  �� ��       ��  h�      ��  h� i       ��  � �!                    �                            � ) * * � - � - � / 0 0 �   2 3 3 � � 5 6 6 � 8 � 8   : ; ; � >   > ?   ? @ @ � � B C C � E � E � G H H � � J K K � � M N N   � P Q Q   � S T T   � V W W � � Y Z Z � � \ ] ] � _ � _ � a b b � � d e e � � g h h � � j k k � m u m o � o r � r s ~ s t t � u u � z � z { { � ~ ~ s  �    � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � * � � ) � � � � � � � � � � � � � � � � � � � � � � � - � � � � � � � � � � 0 � � � � / � � � � � � � � � 8 � � � � � � H � � J 3 5 � 6 � j � � � � � � ; � k � � � e � @ � � B E � � C � K � � � G � _ � Y � � � � � M � P � S � � W � � � � V � r { � � � � � � Z � � � � � � � \ � � � � � ] � � � � � � � a � � d b h  � g � � � � z � � � t m � � � � � � � � � � � � � � � � � � � o             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 